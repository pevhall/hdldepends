package misc_package;
        // Package contents (parameters, types, tasks, functions)
endpackage
