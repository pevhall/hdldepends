
package del_pkg is 
  constant TEST : natural := 2;
end package;
